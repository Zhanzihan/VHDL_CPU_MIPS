library  ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;

entity cmemory is
port
(
    next_addr_in:in std_logic_vector(7 downto 0);
    cm_data_out:out std_logic_vector(32 downto 0)
);
end cmemory;

architecture Behavioral of cmemory is

begin
    process(next_addr_in)
    begin
        case next_addr_in is
            when X"00" =>
                cm_data_out<="000000000000000000000000000000000000000111110000000001000";
            --fetch
            when X"01" =>
                cm_data_out<=B"00_010_000_000000000_0_0000_00_1_000000_000000_0011111_0_1_00000010_000";
            when X"02"=>
                cm_data_out<=B"01_000_001_000000000_0_0000_00_1_000000_000000_0011111_0_1_00000011_000";
            when X"03"=>
                cm_data_out<=B"00_000_000_000000000_1_0000_00_1_000000_000000_0011111_0_1_00000100_000";
            when X"04"=>
                cm_data_out<=B"00_000_000_000000000_0_0000_00_0_000000_000000_0011111_0_0_00000000_100";
            --间址
            when X"05"=>
                cm_data_out<=B"00_100_000_000000000_0_0000_00_1_000000_000000_0011111_0_1_00000101_000";
            when X"06"=>
                cm_data_out<=B"01_000_000_000000000_0_0000_00_1_000000_000000_0011111_0_1_00000110_000";
            when X"07"=>
                cm_data_out<=B"00_001_000_000000000_0_0000_00_1_000000_000000_0011111_0_0_00000000_001";
            --中断
            when X"08"=>    
            when X"09"=>   
            --addu
            when X"0a"=>
                cm_data_out<=B"00_000_000_000000000_0_0000_00_1_100000_100000_1000000_0_0_00000001_010";
            --ori
            when X"0b"=>
                cm_data_out<=B"00_000_000_000000000_0_0111_10_1_100000_000000_0100000_0_0_00000001_010";
            --bne
            when X"0c"=>
                cm_data_out<=B"11_000_000_000000000_0_1110_10_1_000000_000000_0000001_0_0_00001101_000";
            when X"0d"=>
                cm_data_out<=B"10_000_000_000000000_0_0000_00_0_000000_000000_0011111_0_0_00001110_000";
            when X"0e"=>
                cm_data_out<=B"11_000_000_000000000_0_0000_01_1_000001_000000_0000001_0_0_00001111_000";
            when X"0f"=>
                cm_data_out<=B"00_000_000_000000000_1_0100_00_1_100000_100000_0011111_0_0_00010000_000";
            when X"10"=>
                cm_data_out<=B"00_000_000_000000010_0_0000_00_0_000000_000000_0011111_0_0_00011000_000";
            --lw
            when X"11"=>
                cm_data_out<=B"00_011_000_000000000_0_0000_10_0_100000_000000_0011111_0_1_00010010_000";
            when X"12"=>
                cm_data_out<=B"01_000_000_000000000_0_0000_00_0_000000_000000_0011111_0_1_00010011_000";
            when X"13"=>
                cm_data_out<=B"00_000_000_000000000_0_0000_00_0_000000_000000_0100000_0_0_00000001_010";

            --sw
            when X"14"=>
                cm_data_out<=B"00_011_000_000000000_0_0000_10_0_100000_000000_0011111_0_0_00010101_000";
                
            when X"15"=>
                cm_data_out<=B"11_000_000_000000000_0_1110_00_0_000000_100000_0011111_0_0_00010110_000";
            when X"16"=>
                cm_data_out<=B"00_000_000_000000000_0_0000_00_0_000000_000000_0011111_1_0_00000001_010";
            
            --lui
            when X"17"=>
                cm_data_out<=B"00_000_000_000000000_0_1111_10_1_000000_100000_0100000_0_0_00000001_010";
            
            when X"18"=>
                cm_data_out<=B"00_000_000_000000000_0_0000_00_0_000000_000000_0011111_0_0_00000001_010";
            
            when others=>
                cm_data_out<="000000000000000000000000000000000000000111110000000001000";

            end case;
    end process;

end Behavioral;