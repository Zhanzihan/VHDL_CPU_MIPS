library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity overflowReg is
    port (
        
    );
end entity overflowReg;

architecture rtl of overflowReg is
    
begin
    
    
    
end architecture rtl;